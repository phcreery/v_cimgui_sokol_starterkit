module glue

import sokol.gfx

fn C.sapp_sgcontext() gfx.ContextDesc
