module sokolext

import libs.sokolext.c

const (
	imgui_used_import = c.used_import
)
