module sokolext

import libs.sokolext.c as _
